** Profile: "SCHEMATIC1-Parametric"  [ D:\University Projects\OrCAD Projects\Final-Schmitt-Trigger\schmitt-trigger-pspicefiles\schematic1\parametric.sim ] 

** Creating circuit file "Parametric.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3ms 0 SKIPBP 
.STEP LIN PARAM SET 0 1 0.2 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END

** Profile: "SCHEMATIC1-Worst-Case"  [ D:\University Projects\OrCAD Projects\Final-Schmitt-Trigger\Schmitt-Trigger-PSpiceFiles\SCHEMATIC1\Worst-Case.sim ] 

** Creating circuit file "Worst-Case.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3ms 0 SKIPBP 
.WCASE TRAN V([OUT]) YMAX VARY BOTH  HI 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
